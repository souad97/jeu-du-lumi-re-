library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
 
ENTITY LED IS
PORT(
CLOCK_50: IN STD_LOGIC;
LEDG: OUT STD_LOGIC_VECTOR(7 downto 0);
LEDR:OUT STD_LOGIC_VECTOR(9 downto 0);
KEY:IN STD_LOGIC_VECTOR(3 downto 0)
);
 
END LED;
 
 
ARCHITECTURE COUNTER OF LED IS
SIGNAL PRESCALER : INTEGER RANGE 0 TO 500000:=0;
SIGNAL RESULT: INTEGER RANGE 0 TO 1023:=0;
BEGIN
 
PROCESS(CLOCK_50)
BEGIN
IF(CLOCK_50'EVENT AND CLOCK_50='1')THEN
  IF(PRESCALER<500000)THEN
	  PRESCALER<=PRESCALER+1;
	  ELSE
	  PRESCALER<=0;
  END IF;
  IF(PRESCALER=0)THEN
 
     CASE KEY(0) IS
	   WHEN '0' =>
			IF(RESULT<1023)THEN
			 RESULT<=RESULT+1;
			ELSE
			 RESULT<=0;
			END IF;
		WHEN '1'=>
			IF(RESULT>0)THEN
			 RESULT<=RESULT-1;
			ELSE
			 RESULT<=1023;
			END IF;
	  END CASE;
  END IF;
 
END IF;
END PROCESS;
 
PROCESS(CLOCK_50)
BEGIN
IF(CLOCK_50'EVENT AND CLOCK_50='1')THEN
   IF(KEY(1)='0')THEN
	LEDR<= STD_LOGIC_VECTOR(to_unsigned(RESULT,10));
	ELSE
	 FOR i IN 1 TO 10 LOOP
	   IF(RESULT>102*i)THEN
			LEDR(i-1)<='1';
			ELSE
			LEDR(i-1)<='0';
	   END IF;
	 END LOOP;
 
	END IF;
 
 
END IF;
 
 
 
 
 
END PROCESS;
END COUNTER;
